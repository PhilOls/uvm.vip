//
// Template for UVM-compliant interface
//

`ifndef base_if__SV
`define base_if__SV

interface base_if ();

endinterface

`endif
